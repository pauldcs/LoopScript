CLICK
	(540, 240)
	(540, 240)
	(1.0, 1.5);

WRITE
	"hello world";

WAIT	3;

WRITE_RSTR 20;

WRITE_RTEXT 4;